bind CPUtop SIMD_assertions sva_bind (clk, rst, instruction_in, data_in, data_out, instruction_address, data_address, data_R, data_W, done, opcode, CMD_addition, CMD_substruction, CMD_multiplication, CMD_mul_accumulation, CMD_logic_shift_left, CMD_logic_shift_right, CMD_and, CMD_or, CMD_not, CMD_loopjump, CMD_setloop, CMD_load, CMD_store, CMD_set, current_state, STATE_IDLE, STATE_IF, STATE_ID, STATE_EX, STATE_MEM, STATE_HALT, rdata_en, wdata_en);
